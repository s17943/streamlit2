���:      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.2.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��	RestingBP��Cholesterol��MaxHR��Oldpeak�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh&hNhJ�
hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h4�f8�����R�(KhKNNNJ����J����K t�b�C              �?�t�bhOh(�scalar���hJC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hK�
node_count�K�nodes�h*h-K ��h/��R�(KK��h4�V56�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h{hJK ��h|hJK��h}hJK��h~h[K��hh[K ��h�hJK(��h�h[K0��uK8KKt�b�BH                            @E@j8je3�?�           ��@                          �?P>�7���?L            @]@                           @O@d}h���?             E@������������������������       �r�q��?             B@������������������������       �      �?             @                           c@H0sE�d�?0            �R@������������������������       �      �?(             P@������������������������       ����|���?             &@	                        pff�?�ؗ���?�           H�@
                          �}@�@o-4�?�            �s@������������������������       �~�Kƛj�?�            0s@������������������������       �                     @                          �b@^T�7���?�            s@������������������������       ��������?�            @n@������������������������       ��G��l��?'            �O@�t�b�values�h*h-K ��h/��R�(KKKK��h[�C�     Ps@     �z@      1@      Y@      "@     �@@      @      >@      @      @       @     �P@      @      N@      @      @     @r@     Pt@      m@     �S@      m@     �R@              @     �M@     �n@      :@      k@     �@@      >@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ/��hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                            �`@4�5����?�           ��@                          �f@�������?�            �s@                           `@      �?E             Z@������������������������       ��:nR&y�??            �W@������������������������       ��q�q�?             "@                          `[@
Y�+ߧ�?�            �j@������������������������       ���hJ,�?)             Q@������������������������       �&���7��?c            `b@	                        ����?l�?���?�            �y@
                          @g@V��T���?�            �p@������������������������       �F.< ?�?�            �p@������������������������       �                     @                          s@^H���+�?]            �b@������������������������       ����qK�?U            �`@������������������������       �������?             .@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�     �t@     y@     @Q@     @o@      *@     �V@      @      V@      @      @      L@     �c@      $@      M@      G@     @Y@     �p@     �b@     �j@     �K@     �j@      J@              @      J@      X@     �D@      W@      &@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJu�7hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                            �`@p�Vv���?�           ��@                        ����?�dG��?�            �t@                           �I@�ݜ����?M            �]@������������������������       ��q�q�?            �F@������������������������       �z�7�Z�?3            @R@                          P`@�����?�            `j@������������������������       ���f��??            @V@������������������������       � @|���?P            �^@	                           @L@���Q��?           Py@
                          �c@4;����?�            �p@������������������������       ���C���?`            �a@������������������������       �^f�(�7�?M            @_@                        ����?�)z� ��?V            `a@������������������������       �^n����?&             N@������������������������       �p`q�q��?0            �S@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�     @t@     �y@     @T@      o@      L@      O@      >@      .@      :@     �G@      9@     @g@      2@     �Q@      @     �\@     `n@     @d@     @g@      T@      U@     �L@     �Y@      7@     �L@     �T@     �D@      3@      0@     �O@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ��!XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                          ����?U�ք�?�           ��@                          `_@��R�{�?�             w@                          Pe@"Ae���?A            �W@������������������������       ����}<S�?             G@������������������������       ��q�q�?%             H@                          �d@�{WR�&�?�             q@������������������������       ��b��-8�?z            �g@������������������������       ��t����?:            @U@	                           @K@��@�yC�?�            �v@
                          0d@�)O���?Y            �`@������������������������       � 7���B�?             ;@������������������������       �*��ZE�?E            �Z@                           `R@t0�J��?�             m@������������������������       �d�X^_�?�            �l@������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      t@     �y@     �n@     �^@      @@      O@      @      E@      <@      4@     �j@     �N@     @a@     �I@     �R@      $@     @S@     r@      G@     �U@      �?      :@     �F@     �N@      ?@     @i@      <@     @i@      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJC�NhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                          ����?4�5����?�           ��@                          `_@�Ff��K�?�            x@                          `f@�kwY���?G            @Z@������������������������       �r�qG�?D             X@������������������������       �                     "@                        ����?4և����?�            �q@������������������������       �&��ĕu�?�            �n@������������������������       ��ʻ����?             A@	                          �`@�?ʵ���?�            �u@
                          �b@���U��?z            @g@������������������������       �d}h���?_            �a@������������������������       �\X��t�?             G@                          �b@D���\�?p            `d@������������������������       �@4և���?\            �a@������������������������       ��û��|�?             7@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�     �t@     y@      p@     �_@     �E@      O@      A@      O@      "@             �j@     @P@      i@      G@      .@      3@     �R@      q@      L@     @`@      >@     �[@      :@      4@      3@      b@      $@     @`@      "@      ,@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�R�[hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                          ����?6������?�           ��@                          @E@��_���?�             w@                          �c@�S����?$            �L@������������������������       ���k=.��?            �G@������������������������       �                     $@                           @L@�W�o���?�            ps@������������������������       �b�����?�            �k@������������������������       �r�����?;            @V@	                          �`@xƅd�?�            �v@
                          �z@ܷ��?��?~            `i@������������������������       ��j�zZ��?}             i@������������������������       �                      @                          f@噼:��?d            `d@������������������������       �p�ݯ��?]             c@������������������������       �"pc�
�?             &@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�     �t@     �x@      o@     �]@      "@      H@      "@      C@              $@      n@     �Q@     `g@     �A@     �J@      B@     �U@     �q@      5@     �f@      3@     �f@       @             @P@     �X@      L@      X@      "@       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�v}hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                            �^@U�ք�?�           ��@                          �U@����l��?W             a@������������������������       �                     @                          �]@t�U����?V            �`@������������������������       ���?^�k�?)            �Q@������������������������       �     ��?-             P@       
                   �`@h��b#��?v           ��@       	                 ����?02�U;q�?�            �u@������������������������       ��ګH9�?�            �j@������������������������       �<��¤�?Q             a@                          0`@�pX���?�             o@������������������������       �����?D            @[@������������������������       �sYi9��?T            `a@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      t@     �y@      3@     �]@      @              0@     �]@       @      Q@      ,@      I@     �r@     `r@     �j@      a@     �c@      K@      K@     �T@     �V@     �c@      1@      W@     @R@     �P@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJg}�XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                            P`@0����?�           ��@                          �b@�<ݚ�?�            �s@                           `@��8��)�?>            �W@������������������������       ���S�ۿ?;            �V@������������������������       �      �?             @                          �d@X��8��?�            �k@������������������������       �                     @������������������������       �~�1u���?�            @k@	                           @L@�"�,��?	           0z@
                          @E@(הn��?�            �q@������������������������       ����}<S�?             7@������������������������       ��GN�z�?�            �p@                        pff�?�eP*L��?T            �`@������������������������       �^����?            �E@������������������������       ��VM�?9            @V@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      u@     �x@     �Q@     �n@      "@     @U@      @      U@      @      �?     �N@      d@      @              M@      d@     �p@      c@     �i@     @T@       @      5@     �i@      N@      N@      R@      ?@      (@      =@      N@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ	�tlhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                          ����?�+	G�?�           ��@                          `_@�ɞ`s�?�            �v@                            J@r�����?9            @V@������������������������       ���}*_��?             ;@������������������������       �V��z4�?)             O@                          @E@�I;F���?�            Pq@������������������������       �        
             3@������������������������       ��T|n�q�?�             p@	                          �b@2�K36��?�             w@
                           �R@h8"J{�?�            �r@������������������������       ��X�3�m�?�            pr@������������������������       ��q�q�?             @                          0c@��
P��?)            �Q@������������������������       �                      @������������������������       �`՟�G��?$             O@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�     `t@     �y@     �o@     �\@      B@     �J@      1@      $@      3@     �E@      k@     �N@              3@      k@      E@     �R@     `r@      C@     @p@      B@     0p@       @      �?      B@      A@       @              <@      A@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�ޡhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                             @L@6������?�           ��@                        ����?h�����?&            |@                          �Z@ά��.��?�            @p@������������������������       �����X�?	             ,@������������������������       �"�W1��?�            �n@                          @e@V��N��?�            �g@������������������������       ���p\�?            �D@������������������������       ������?g            `b@	                        ����?��
n��?�            �q@
                          �`@)O���?E             [@������������������������       ��GN�z�?             6@������������������������       ��&!��?6            �U@                          �s@d��o�t�?u            @f@������������������������       �,���i�?m            �d@������������������������       �X�Cc�?             ,@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�     �t@     �x@      o@     �h@     �h@     �N@      @      $@     `h@     �I@      I@     @a@      @      C@     �G@      Y@     �U@      i@     �L@     �I@      @      1@      J@      A@      =@     �b@      4@      b@      "@      @�t�bubhhubehhub.